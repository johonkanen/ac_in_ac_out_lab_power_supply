LIBRARY ieee  ; 
    USE ieee.NUMERIC_STD.all  ; 
    USE ieee.std_logic_1164.all  ; 
    use ieee.math_real.all;

package buck_sw_model_pkg is

end package;

package body buck_sw_model_pkg is

end package body;
